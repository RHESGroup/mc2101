--This file is automatically generated, please do not change the content
--file content description:
--boot code for flash
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
PACKAGE CONSTANTS IS
TYPE c_mem IS ARRAY (0 TO 2**12 -1) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
CONSTANT boot_code : c_mem:=(
x"6F",
x"00",
x"80",
x"30",
x"6F",
x"00",
x"80",
x"47",
x"6F",
x"00",
x"80",
x"4A",
x"6F",
x"00",
x"40",
x"47",
x"6F",
x"00",
x"00",
x"4A",
x"6F",
x"00",
x"C0",
x"49",
x"6F",
x"00",
x"80",
x"49",
x"6F",
x"00",
x"40",
x"49",
x"6F",
x"00",
x"00",
x"49",
x"6F",
x"00",
x"00",
x"46",
x"6F",
x"00",
x"80",
x"48",
x"6F",
x"00",
x"40",
x"48",
x"6F",
x"00",
x"00",
x"48",
x"6F",
x"00",
x"C0",
x"47",
x"6F",
x"00",
x"80",
x"47",
x"6F",
x"00",
x"40",
x"47",
x"6F",
x"00",
x"00",
x"47",
x"6F",
x"00",
x"C0",
x"46",
x"6F",
x"00",
x"80",
x"46",
x"6F",
x"00",
x"40",
x"46",
x"6F",
x"00",
x"00",
x"46",
x"6F",
x"00",
x"C0",
x"45",
x"6F",
x"00",
x"80",
x"45",
x"6F",
x"00",
x"40",
x"45",
x"6F",
x"00",
x"00",
x"45",
x"6F",
x"00",
x"C0",
x"44",
x"6F",
x"00",
x"80",
x"44",
x"6F",
x"00",
x"40",
x"44",
x"6F",
x"00",
x"00",
x"44",
x"6F",
x"00",
x"C0",
x"43",
x"6F",
x"00",
x"80",
x"43",
x"6F",
x"00",
x"40",
x"43",
x"6F",
x"00",
x"00",
x"43",
x"6F",
x"00",
x"C0",
x"42",
x"6F",
x"00",
x"80",
x"42",
x"6F",
x"00",
x"40",
x"42",
x"6F",
x"00",
x"00",
x"42",
x"6F",
x"00",
x"C0",
x"41",
x"6F",
x"00",
x"80",
x"41",
x"6F",
x"00",
x"40",
x"41",
x"6F",
x"00",
x"00",
x"41",
x"6F",
x"00",
x"C0",
x"40",
x"6F",
x"00",
x"80",
x"40",
x"6F",
x"00",
x"40",
x"40",
x"6F",
x"00",
x"00",
x"40",
x"6F",
x"00",
x"C0",
x"3F",
x"6F",
x"00",
x"80",
x"3F",
x"6F",
x"00",
x"40",
x"3F",
x"6F",
x"00",
x"00",
x"3F",
x"6F",
x"00",
x"C0",
x"3D",
x"6F",
x"00",
x"80",
x"3D",
x"6F",
x"00",
x"40",
x"3D",
x"6F",
x"00",
x"00",
x"3D",
x"6F",
x"00",
x"C0",
x"3C",
x"6F",
x"00",
x"80",
x"3C",
x"6F",
x"00",
x"40",
x"3C",
x"6F",
x"00",
x"00",
x"3C",
x"6F",
x"00",
x"C0",
x"3B",
x"6F",
x"00",
x"80",
x"3B",
x"6F",
x"00",
x"40",
x"3B",
x"6F",
x"00",
x"00",
x"3B",
x"6F",
x"00",
x"C0",
x"3A",
x"6F",
x"00",
x"80",
x"3A",
x"6F",
x"00",
x"40",
x"3A",
x"6F",
x"00",
x"00",
x"3A",
x"B7",
x"00",
x"10",
x"00",
x"13",
x"01",
x"10",
x"00",
x"23",
x"A0",
x"20",
x"00",
x"13",
x"01",
x"00",
x"00",
x"03",
x"A1",
x"00",
x"00",
x"93",
x"01",
x"11",
x"00",
x"23",
x"A0",
x"30",
x"00",
x"93",
x"01",
x"00",
x"00",
x"83",
x"A1",
x"00",
x"00",
x"13",
x"82",
x"11",
x"00",
x"23",
x"A0",
x"40",
x"00",
x"13",
x"02",
x"00",
x"00",
x"03",
x"A2",
x"00",
x"00",
x"93",
x"02",
x"12",
x"00",
x"23",
x"A0",
x"50",
x"00",
x"93",
x"02",
x"00",
x"00",
x"83",
x"A2",
x"00",
x"00",
x"13",
x"83",
x"12",
x"00",
x"23",
x"A0",
x"60",
x"00",
x"13",
x"03",
x"00",
x"00",
x"03",
x"A3",
x"00",
x"00",
x"93",
x"03",
x"13",
x"00",
x"23",
x"A0",
x"70",
x"00",
x"93",
x"03",
x"00",
x"00",
x"83",
x"A3",
x"00",
x"00",
x"13",
x"84",
x"13",
x"00",
x"23",
x"A0",
x"80",
x"00",
x"13",
x"04",
x"00",
x"00",
x"03",
x"A4",
x"00",
x"00",
x"93",
x"04",
x"14",
x"00",
x"23",
x"A0",
x"90",
x"00",
x"93",
x"04",
x"00",
x"00",
x"83",
x"A4",
x"00",
x"00",
x"13",
x"85",
x"14",
x"00",
x"23",
x"A0",
x"A0",
x"00",
x"13",
x"05",
x"00",
x"00",
x"03",
x"A5",
x"00",
x"00",
x"93",
x"05",
x"15",
x"00",
x"23",
x"A0",
x"B0",
x"00",
x"93",
x"05",
x"00",
x"00",
x"83",
x"A5",
x"00",
x"00",
x"13",
x"86",
x"15",
x"00",
x"23",
x"A0",
x"C0",
x"00",
x"13",
x"06",
x"00",
x"00",
x"03",
x"A6",
x"00",
x"00",
x"93",
x"06",
x"16",
x"00",
x"23",
x"A0",
x"D0",
x"00",
x"93",
x"06",
x"00",
x"00",
x"83",
x"A6",
x"00",
x"00",
x"13",
x"87",
x"16",
x"00",
x"23",
x"A0",
x"E0",
x"00",
x"13",
x"07",
x"00",
x"00",
x"03",
x"A7",
x"00",
x"00",
x"93",
x"07",
x"17",
x"00",
x"23",
x"A0",
x"F0",
x"00",
x"93",
x"07",
x"00",
x"00",
x"83",
x"A7",
x"00",
x"00",
x"13",
x"88",
x"17",
x"00",
x"23",
x"A0",
x"00",
x"01",
x"13",
x"08",
x"00",
x"00",
x"03",
x"A8",
x"00",
x"00",
x"93",
x"08",
x"18",
x"00",
x"23",
x"A0",
x"10",
x"01",
x"93",
x"08",
x"00",
x"00",
x"83",
x"A8",
x"00",
x"00",
x"13",
x"89",
x"18",
x"00",
x"23",
x"A0",
x"20",
x"01",
x"13",
x"09",
x"00",
x"00",
x"03",
x"A9",
x"00",
x"00",
x"93",
x"09",
x"19",
x"00",
x"23",
x"A0",
x"30",
x"01",
x"93",
x"09",
x"00",
x"00",
x"83",
x"A9",
x"00",
x"00",
x"13",
x"8A",
x"19",
x"00",
x"23",
x"A0",
x"40",
x"01",
x"13",
x"0A",
x"00",
x"00",
x"03",
x"AA",
x"00",
x"00",
x"93",
x"0A",
x"1A",
x"00",
x"23",
x"A0",
x"50",
x"01",
x"93",
x"0A",
x"00",
x"00",
x"83",
x"AA",
x"00",
x"00",
x"13",
x"8B",
x"1A",
x"00",
x"23",
x"A0",
x"60",
x"01",
x"13",
x"0B",
x"00",
x"00",
x"03",
x"AB",
x"00",
x"00",
x"93",
x"0B",
x"1B",
x"00",
x"23",
x"A0",
x"70",
x"01",
x"93",
x"0B",
x"00",
x"00",
x"83",
x"AB",
x"00",
x"00",
x"13",
x"8C",
x"1B",
x"00",
x"23",
x"A0",
x"80",
x"01",
x"13",
x"0C",
x"00",
x"00",
x"03",
x"AC",
x"00",
x"00",
x"93",
x"0C",
x"1C",
x"00",
x"23",
x"A0",
x"90",
x"01",
x"93",
x"0C",
x"00",
x"00",
x"83",
x"AC",
x"00",
x"00",
x"13",
x"8D",
x"1C",
x"00",
x"23",
x"A0",
x"A0",
x"01",
x"13",
x"0D",
x"00",
x"00",
x"03",
x"AD",
x"00",
x"00",
x"93",
x"0D",
x"1D",
x"00",
x"23",
x"A0",
x"B0",
x"01",
x"93",
x"0D",
x"00",
x"00",
x"83",
x"AD",
x"00",
x"00",
x"13",
x"8E",
x"1D",
x"00",
x"23",
x"A0",
x"C0",
x"01",
x"13",
x"0E",
x"00",
x"00",
x"03",
x"AE",
x"00",
x"00",
x"93",
x"0E",
x"1E",
x"00",
x"23",
x"A0",
x"D0",
x"01",
x"93",
x"0E",
x"00",
x"00",
x"83",
x"AE",
x"00",
x"00",
x"13",
x"8F",
x"1E",
x"00",
x"23",
x"A0",
x"E0",
x"01",
x"13",
x"0F",
x"00",
x"00",
x"03",
x"AF",
x"00",
x"00",
x"93",
x"0F",
x"1F",
x"00",
x"23",
x"A0",
x"F0",
x"01",
x"93",
x"0F",
x"00",
x"00",
x"83",
x"AF",
x"00",
x"00",
x"93",
x"0F",
x"20",
x"01",
x"23",
x"80",
x"F0",
x"01",
x"93",
x"0F",
x"00",
x"01",
x"83",
x"8F",
x"00",
x"00",
x"23",
x"90",
x"F0",
x"01",
x"93",
x"8F",
x"0F",
x"00",
x"83",
x"9F",
x"00",
x"00",
x"6F",
x"00",
x"00",
x"00",
x"93",
x"00",
x"00",
x"18",
x"93",
x"90",
x"40",
x"00",
x"F3",
x"90",
x"00",
x"30",
x"F3",
x"D0",
x"58",
x"30",
x"93",
x"00",
x"00",
x"00",
x"13",
x"81",
x"00",
x"00",
x"93",
x"81",
x"00",
x"00",
x"13",
x"82",
x"00",
x"00",
x"93",
x"82",
x"00",
x"00",
x"13",
x"83",
x"00",
x"00",
x"93",
x"83",
x"00",
x"00",
x"13",
x"84",
x"00",
x"00",
x"93",
x"84",
x"00",
x"00",
x"13",
x"85",
x"00",
x"00",
x"93",
x"85",
x"00",
x"00",
x"13",
x"86",
x"00",
x"00",
x"93",
x"86",
x"00",
x"00",
x"13",
x"87",
x"00",
x"00",
x"93",
x"87",
x"00",
x"00",
x"13",
x"88",
x"00",
x"00",
x"93",
x"88",
x"00",
x"00",
x"13",
x"89",
x"00",
x"00",
x"93",
x"89",
x"00",
x"00",
x"13",
x"8A",
x"00",
x"00",
x"93",
x"8A",
x"00",
x"00",
x"13",
x"8B",
x"00",
x"00",
x"93",
x"8B",
x"00",
x"00",
x"13",
x"8C",
x"00",
x"00",
x"93",
x"8C",
x"00",
x"00",
x"13",
x"8D",
x"00",
x"00",
x"93",
x"8D",
x"00",
x"00",
x"13",
x"8E",
x"00",
x"00",
x"93",
x"8E",
x"00",
x"00",
x"13",
x"8F",
x"00",
x"00",
x"93",
x"8F",
x"00",
x"00",
x"17",
x"11",
x"10",
x"00",
x"13",
x"01",
x"C1",
x"C6",
x"17",
x"0D",
x"10",
x"00",
x"13",
x"0D",
x"4D",
x"C6",
x"97",
x"0D",
x"10",
x"00",
x"93",
x"8D",
x"CD",
x"C5",
x"63",
x"58",
x"BD",
x"01",
x"23",
x"20",
x"0D",
x"00",
x"13",
x"0D",
x"4D",
x"00",
x"E3",
x"DC",
x"AD",
x"FF",
x"13",
x"05",
x"00",
x"00",
x"93",
x"05",
x"00",
x"00",
x"93",
x"03",
x"00",
x"00",
x"B7",
x"03",
x"FF",
x"FF",
x"F3",
x"A3",
x"43",
x"30",
x"93",
x"03",
x"80",
x"00",
x"F3",
x"A3",
x"03",
x"30",
x"93",
x"03",
x"00",
x"00",
x"EF",
x"F0",
x"9F",
x"D2",
x"6F",
x"00",
x"00",
x"00",
x"23",
x"20",
x"31",
x"00",
x"23",
x"22",
x"41",
x"00",
x"23",
x"24",
x"51",
x"00",
x"23",
x"26",
x"61",
x"00",
x"23",
x"28",
x"71",
x"00",
x"23",
x"2A",
x"A1",
x"00",
x"23",
x"2C",
x"B1",
x"00",
x"23",
x"2E",
x"C1",
x"00",
x"23",
x"20",
x"D1",
x"02",
x"23",
x"22",
x"E1",
x"02",
x"23",
x"24",
x"F1",
x"02",
x"23",
x"26",
x"01",
x"03",
x"23",
x"28",
x"11",
x"03",
x"23",
x"2A",
x"C1",
x"03",
x"23",
x"2C",
x"D1",
x"03",
x"23",
x"2E",
x"E1",
x"03",
x"23",
x"20",
x"F1",
x"05",
x"67",
x"80",
x"00",
x"00",
x"83",
x"21",
x"01",
x"00",
x"03",
x"22",
x"41",
x"00",
x"83",
x"22",
x"81",
x"00",
x"03",
x"23",
x"C1",
x"00",
x"83",
x"23",
x"01",
x"01",
x"03",
x"25",
x"41",
x"01",
x"83",
x"25",
x"81",
x"01",
x"03",
x"26",
x"C1",
x"01",
x"83",
x"26",
x"01",
x"02",
x"03",
x"27",
x"41",
x"02",
x"83",
x"27",
x"81",
x"02",
x"03",
x"28",
x"C1",
x"02",
x"83",
x"28",
x"01",
x"03",
x"03",
x"2E",
x"41",
x"03",
x"83",
x"2E",
x"81",
x"03",
x"03",
x"2F",
x"C1",
x"03",
x"83",
x"2F",
x"01",
x"04",
x"83",
x"20",
x"41",
x"04",
x"13",
x"01",
x"81",
x"04",
x"73",
x"00",
x"20",
x"30",
x"6F",
x"00",
x"00",
x"00",
x"6F",
x"00",
x"00",
x"00",
x"13",
x"01",
x"81",
x"FB",
x"23",
x"22",
x"11",
x"04",
x"EF",
x"F0",
x"9F",
x"F5",
x"F3",
x"63",
x"10",
x"34",
x"93",
x"83",
x"43",
x"00",
x"F3",
x"93",
x"13",
x"34",
x"6F",
x"F0",
x"1F",
x"F9",
x"13",
x"01",
x"81",
x"FB",
x"23",
x"22",
x"11",
x"04",
x"EF",
x"F0",
x"DF",
x"F3",
x"6F",
x"F0",
x"1F",
x"F8",
x"6F",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00");
END PACKAGE CONSTANTS;
